module and_design( a, b, c);
input a,b;
output c;
assign c=a&b;
endmodule:and_design

