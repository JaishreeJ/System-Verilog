module top();
and_if inf();
and_design a1 (.a(inf.a),.b(inf.b),.c(inf.c));
tb_and a2 (inf);
endmodule:top
