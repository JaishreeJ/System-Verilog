module modport_design(mod_intr inf);
assign inf.dut.c=(inf.dut.a)&(inf.dut.b);
endmodule:modport_design


