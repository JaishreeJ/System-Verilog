module modport_top();
mod_intr inf();
modport_design a1(inf);
modport_tb a2(inf);
endmodule:modport_top

