
interface and_if;
logic a,b;
logic c;
endinterface:and_if

