module repeat_for;
initial begin
  for (int i = 1;i<=4;i++)begin   
    $display ("Good morning");   
    $display ("Keep Shining");
  end 
end 
endmodule 

